module or_gate (a,b,y);

input wire a;
input wire b;
output wire y;
assign y = a|b;

endmodule